
module nios (
	clk_clk,
	ps2_loc_export,
	reset_reset_n);	

	input		clk_clk;
	output	[4:0]	ps2_loc_export;
	input		reset_reset_n;
endmodule
